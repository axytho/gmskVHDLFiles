--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   17:58:37 04/21/2020
-- Design Name:   
-- Module Name:   /users/students/r0666113/Documents/gmsk100-digital/xilinx/vhdlGroup4FirstRun/hann_filter_tb.vhd
-- Project Name:  vhdlGroup4FirstRun
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: hann_filter
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
USE ieee.numeric_std.ALL;
 
ENTITY full_simulation_tb IS
END full_simulation_tb;
 
ARCHITECTURE behavior OF full_simulation_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
--    COMPONENT hann_filter
--    PORT(
--         clk : IN  std_logic;
--         inputValue : IN  signed(7 downto 0);
--         newValue : IN  std_logic;
--         outputValue : OUT  signed(7 downto 0);
--         doneFull : OUT  std_logic
--        );
--    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal input_I : signed(7 downto 0) := "00000000";
	signal input_Q : signed(7 downto 0) := "00000000";
   signal newValue : std_logic := '0';
	signal start_atan : std_logic := '0';

 	--Outputs
   signal output_I : signed(7 downto 0);
	signal output_Q : signed(7 downto 0);
   signal done_I : std_logic;
	signal done_Q : std_logic;
	signal done_arctan : std_logic;
	signal angle_out : signed(7 downto 0);
	

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut_I: entity work.low_pass_filter_22 PORT MAP (
          clk => clk,
          inputValue => input_I,
          newValue => newValue,
          outputValue => output_I,
          doneFull => done_I
        );
		  
	 uut_Q: entity work.low_pass_filter_22 PORT MAP (
          clk => clk,
          inputValue => input_Q,
          newValue => newValue,
          outputValue => output_Q,
          doneFull => done_Q
        );

    atan_cordic_uut: entity work.atan_cordic_full_circle port map(
		clk => clk,
		inputXFull => output_I,
		inputYFull => output_Q,
		startFull => start_atan,
		doneFull => done_arctan,
		angleFull => angle_out
	);	  
	
	rising_edge_to_arctan: entity work.rising_edge_block port map(
	    clk => clk,
		 signal_in => done_I,
		 rising_edge_signal => start_atan
	);

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
	
	newValue_process :process
   begin
		newValue <= '0';
		wait for 19990 ns;
		newValue <= '1';
		wait for 10 ns;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;
		--WARNING: stops being accurate after 13 ms (MATLAB time) or 1.3 ms (VHDL time)
		
		input_I <= "00010000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00001101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00001011"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00001010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00001001"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00001000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00001110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000110"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00010000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "00000101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001111"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00001011"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00001101"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00001100"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "00001001"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00001010"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00001000"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000011"; 
 wait for 20000 ns; 
 input_I <= "11110000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "00000110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "00000100"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110001"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110010"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "11110111"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000010"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110101"; 
 input_Q <= "11110101"; 
 wait for 20000 ns; 
 input_I <= "11110111"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "11111010"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111110"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000001"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111100"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111100"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111110"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111011"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111000"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110100"; 
 wait for 20000 ns; 
 input_I <= "11111000"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "11111011"; 
 input_Q <= "11110001"; 
 wait for 20000 ns; 
 input_I <= "11111111"; 
 input_Q <= "11110010"; 
 wait for 20000 ns; 
 input_I <= "00000010"; 
 input_Q <= "11110011"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "00000100"; 
 input_Q <= "11111010"; 
 wait for 20000 ns; 
 input_I <= "00000011"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "00000000"; 
 input_Q <= "00000000"; 
 wait for 20000 ns; 
 input_I <= "11111101"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11111001"; 
 input_Q <= "00000001"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11111111"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11111101"; 
 wait for 20000 ns; 
 input_I <= "11110011"; 
 input_Q <= "11111001"; 
 wait for 20000 ns; 
 input_I <= "11110100"; 
 input_Q <= "11110110"; 
 wait for 20000 ns; 
 input_I <= "11110110"; 
 input_Q <= "11110011"; 
		
		
		
		
 end process;
END;
